`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/07/21 21:47:06
// Design Name: 
// Module Name: spi_transfer
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module spi_transfer(
//	input wire sys_clk,
//	input wire rst_n,
//	input wire [7:0] data,
//	output
//    );
//endmodule
